from https://naif.jpl.nasa.gov/naif/toolkit_FORTRAN.html
